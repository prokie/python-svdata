module ansi_module_a (
  input var logic a,
  input var logic b
);
  
endmodule